//  Class: wdog_ref_model
//
class wdog_ref_model extends uvm_component;
    `uvm_component_utils(wdog_ref_model);

    // TODO: Implementation of ref model
    //  Group: Components


    //  Group: Variables


    //  Group: Functions

    //  Constructor: new
    function new(string name = "wdog_ref_model", uvm_component parent);
        super.new(name, parent);
    endfunction: new

    
endclass: wdog_ref_model
